
module twox1Mux(
  input [31:0] A,B,
  input SEL,
  output reg[31:0] Y);
  always @ (A or B or SEL)
    begin 
      if (SEL==0)
        Y=A;
      else
        Y=B;
    end
endmodule